// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
// Created on Sun Nov 24 14:30:19 2024

// synthesis message_off 10175

`timescale 1ns/1ns

module controller (
    clock,reset,TC,B,
    T3,T9,W,H,R,Y,G);

    input clock;
    input reset;
    input TC;
    input B;
    tri0 reset;
    tri0 TC;
    tri0 B;
    output T3;
    output T9;
    output W;
    output H;
    output R;
    output Y;
    output G;
    reg T3;
    reg T9;
    reg W;
    reg H;
    reg R;
    reg Y;
    reg G;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter yellow=0,red=1,green=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or TC or B)
    begin
        if (reset) begin
            reg_fstate <= green;
            T3 <= 1'b0;
            T9 <= 1'b0;
            W <= 1'b0;
            H <= 1'b0;
            R <= 1'b0;
            Y <= 1'b0;
            G <= 1'b0;
        end
        else begin
            T3 <= 1'b0;
            T9 <= 1'b0;
            W <= 1'b0;
            H <= 1'b0;
            R <= 1'b0;
            Y <= 1'b0;
            G <= 1'b0;
            case (fstate)
                yellow: begin
                    if (TC)
                        reg_fstate <= red;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= yellow;

                    H <= 1'b1;

                    T9 <= TC;

                    Y <= 1'b1;
                end
                red: begin
                    if (TC)
                        reg_fstate <= green;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= red;

                    R <= 1'b1;

                    W <= 1'b1;
                end
                green: begin
                    if (B)
                        reg_fstate <= yellow;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= green;

                    T3 <= B;

                    H <= 1'b1;

                    G <= 1'b1;
                end
                default: begin
                    T3 <= 1'bx;
                    T9 <= 1'bx;
                    W <= 1'bx;
                    H <= 1'bx;
                    R <= 1'bx;
                    Y <= 1'bx;
                    G <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // controller
